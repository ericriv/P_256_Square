

module P_256_Square_tb();

	


	initial begin
	#20 $stop;
	end 

endmodule