

module P_256_Square(

);



endmodule