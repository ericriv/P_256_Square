

module P_256_Square_tb();



endmodule