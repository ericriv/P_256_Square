

module P_256_Reducer(

);

endmodule
